**** Altos spice deck for characterization release 19.1.2.294
***            
*** Info_arc:

.temp 25

V4 5 0 pwl(0 0 1e-10 1.8)
C4 6 0 1.12151e-14
.ic v(6) = 1.8
MXM0.xsky130_fd_pr__nfet_01v8.msky130_fd_pr__nfet_01v8_0x4 6 5 0 0 inverter:XM0:nfet_01v8:xsky130_fd_pr__nfet_01v8:sky130_fd_pr__nfet_01v8:msky130_fd_pr__nfet_01v8:sky130_fd_pr__nfet_01v8__model L=1.5e-07 W=1e-06 NRS=0 NRD=0 SA=0 SB=0 SD=0 NF=1 
.meas tran AltosDeviceCap00000004 INTEG i(V4) from=0 to=1e-10

V8 10 9 pwl(0 0 1e-10 1.8)
C8 0 10 6.37999e-15
.ic v(0) = 0
MXM1.xsky130_fd_pr__pfet_01v8.msky130_fd_pr__pfet_01v8_0x8 0 9 10 10 inverter:XM1:pfet_01v8:xsky130_fd_pr__pfet_01v8:sky130_fd_pr__pfet_01v8:msky130_fd_pr__pfet_01v8:sky130_fd_pr__pfet_01v8__model L=1.5e-07 W=1.6e-06 NRS=0 NRD=0 SA=0 SB=0 SD=0 NF=1 
.meas tran AltosDeviceCap00000008 INTEG i(V8) from=0 to=1e-10

.model inverter:XM0:nfet_01v8:xsky130_fd_pr__nfet_01v8:sky130_fd_pr__nfet_01v8:msky130_fd_pr__nfet_01v8:sky130_fd_pr__nfet_01v8__model.62 nmos level=54 version=4.5 a0=1.5000000e+00 a1=0.0000000e+00
+  a2=4.2385546e-01 acde=4.0000000e-01 acnqsmod=0 af=1.0000000e+00 agidl=0.0000000e+00
+  ags=1.2500000e+00 aigbacc=1.0000000e+00 aigbinv=3.5000000e-01 aigc=4.3000000e-01 aigsd=4.3000000e-01
+  alpha0=1.9079543e-07 alpha1=8.5000000e-01 at=-3.4212579e+05 b0=0.0000000e+00 b1=0.0000000e+00
+  beta0=9.4472679e+00 bgidl=2.3000000e+09 bigbacc=0.0000000e+00 bigbinv=3.0000000e-02 bigc=5.4000000e-02
+  bigsd=5.4000000e-02 binunit=2 bvs=1.1700000e+01 capmod=2 cdsc=0.0000000e+00
+  cdscb=0.0000000e+00 cdscd=2.0520000e-03 cf=1.4067000e-12 cgbo=1.0000000e-13 cgdl=0.0000000e+00
+  cgdo=2.4490680e-10 cgidl=5.0000000e-01 cgsl=0.0000000e+00 cgso=2.4490680e-10 cigbacc=0.0000000e+00
+  cigbinv=6.0000000e-03 cigc=7.5000000e-02 cigsd=7.5000000e-02 cit=0.0000000e+00 cjs=1.3397492e-03
+  cjswgs=2.3823279e-10 cjsws=3.6735420e-11 ckappas=6.0000000e-01 clc=1.0000000e-07 cle=6.0000000e-01
+  delta=1.0000000e-02 diomod=1 dlc=9.8790800e-09 dlcig=0.0000000e+00 dmcg=0.0000000e+00
+  dmcgt=0.0000000e+00 dmdg=0.0000000e+00 drout=5.0332666e-01 dsub=4.5862506e-01 dvt0=0.0000000e+00
+  dvt0w=-3.5800000e+00 dvt1=5.3000000e-01 dvt1w=1.6706000e+06 dvt2=-3.2000000e-02 dvt2w=6.8000000e-02
+  dvtp0=0.0000000e+00 dvtp1=0.0000000e+00 dwb=0.0000000e+00 dwc=0.0000000e+00 dwg=0.0000000e+00
+  ef=8.4000000e-01 egidl=8.0000000e-01 eigbinv=1.1000000e+00 em=4.1000000e+07 epsrox=3.9000000e+00
+  eta0=6.9413878e-04 etab=-4.3998000e-02 eu=1.6700000e+00 fnoimod=1 fprout=0.0000000e+00
+  gbmin=1.0000000e-12 geomod=0 igbmod=0 igcmod=0 ijthsfwd=1.0000000e-01
+  ijthsrev=1.0000000e-01 jss=2.7500000e-03 jsws=6.0000000e-10 k1=9.0707349e-01 k2=-5.0395190e-02
+  k3=2.0000000e+00 k3b=5.4000000e-01 keta=7.4655023e-01 kf=0.0000000e+00 kt1=1.6188553e-01
+  kt1l=0.0000000e+00 kt2=-2.8878939e-02 ku0=-2.7000000e-08 kvsat=2.0000000e-01 kvth0=9.8000000e-09
+  lalpha0=-2.0282093e-14 lambda=0.0000000e+00 lat=4.8290697e-02 lbeta0=5.5534302e-07 lc=5.0000000e-09
+  lint=1.1932000e-08 lintnoi=-1.0000000e-07 lk2=-8.5802911e-09 lketa=-9.4166860e-08 lkt1=-4.8290697e-08
+  lku0=0.0000000e+00 lkvth0=0.0000000e+00 ll=0.0000000e+00 llc=0.0000000e+00 lln=1.0000000e+00
+  llodku0=0.0000000e+00 llodvth=0.0000000e+00 lmax=1.8000000e-07 lmin=1.5000000e-07 lnfactor=-3.8529747e-06
+  lodeta0=1.0000000e+00 lodk2=1.0000000e+00 lp=1.0000000e+00 lpe0=1.0325000e-07 lpeb=-7.0820000e-08
+  lu0=-6.8814244e-11 lua=-4.2978721e-19 lub=2.2496221e-25 luc=7.0427153e-17 lvsat=-6.7143386e-03
+  lvth0=5.3795596e-08 lw=0.0000000e+00 lwc=0.0000000e+00 lwl=0.0000000e+00 lwlc=0.0000000e+00
+  lwn=1.0000000e+00 minv=0.0000000e+00 mjs=4.4000000e-01 mjswgs=8.0000000e-01 mjsws=9.0000000e-04
+  mobmod=0 moin=6.9000000e+00 ndep=1.7000000e+17 nfactor=3.1183538e+01 ngate=1.0000000e+23
+  ngcon=1.0000000e+00 nigbacc=0.0000000e+00 nigbinv=0.0000000e+00 nigc=0.0000000e+00 njs=1.2928000e+00
+  noff=3.4037000e+00 noia=2.5000000e+42 noib=0.0000000e+00 noic=0.0000000e+00 nsd=1.0000000e+20
+  ntnoi=1.0000000e+00 ntox=1.0000000e+00 palpha0=2.4668745e-20 pat=-5.8735106e-08 pbeta0=-6.7545372e-13
+  pbs=7.2900000e-01 pbswgs=9.5578000e-01 pbsws=2.0000000e-01 pclm=1.8242793e-01 pdiblc1=3.5697215e-01
+  pdiblc2=8.4061121e-03 pdiblcb=-1.0329577e-01 pdits=0.0000000e+00 pditsd=0.0000000e+00 pditsl=0.0000000e+00
+  permod=1 phin=0.0000000e+00 pigcd=1.0000000e+00 pk2=1.0436054e-14 pketa=1.1453346e-13
+  pkt1=5.8735106e-14 pku0=0.0000000e+00 pkvth0=0.0000000e+00 pnfactor=4.6863038e-12 poxedge=1.0000000e+00
+  prt=0.0000000e+00 prwb=0.0000000e+00 prwg=2.1507000e-02 pscbe1=7.9141988e+08 pscbe2=1.0000000e-12
+  pu0=8.3697526e-17 pua=5.2274244e-25 pub=-2.7361749e-31 puc=-8.5659279e-23 pvag=0.0000000e+00
+  pvsat=8.1665291e-09 pvth0=-6.5430615e-14 rbdb=5.0000000e+01 rbodymod=1 rbpb=5.0000000e+01
+  rbpd=5.0000000e+01 rbps=5.0000000e+01 rbsb=5.0000000e+01 rdsmod=0 rdsw=6.5968000e+01
+  rdswmin=0.0000000e+00 rdw=0.0000000e+00 rdwmin=0.0000000e+00 rgatemod=0 rnoia=9.4000000e-01
+  rnoib=2.6000000e-01 rsh=1.0000000e+00 rshg=1.0000000e-01 rsw=0.0000000e+00 rswmin=0.0000000e+00
+  saref=1.0400000e-06 sbref=1.0400000e-06 steta0=0.0000000e+00 stk2=0.0000000e+00 tcj=7.9200000e-04
+  tcjsw=1.0000000e-05 tcjswg=0.0000000e+00 tempmod=0 tku0=0.0000000e+00 tnoia=1.5000000e+07
+  tnoib=9.9000000e+06 tnoimod=1 tnom=3.0000000e+01 toxe=4.1480000e-09 toxm=4.1480000e-09
+  toxref=4.1480000e-09 tpb=1.2287000e-03 tpbsw=0.0000000e+00 tpbswg=0.0000000e+00 trnqsmod=0
+  tvfbsdoff=0.0000000e+00 tvoff=0.0000000e+00 u0=2.8796080e-02 ua=-1.1788768e-09 ua1=-2.3847336e-11
+  ub=1.1212913e-18 ub1=7.0775317e-19 uc=-4.7732100e-10 uc1=1.4718625e-10 ud=0.0000000e+00
+  up=0.0000000e+00 ute=-1.3190432e+00 vbm=-3.0000000e+00 vfbcv=-1.0000000e+00 vfbsdoff=0.0000000e+00
+  voff=-2.0753000e-01 voffcv=-1.7287000e-01 voffl=5.8197729e-09 vsat=2.1519870e+05 vth0=3.1881430e-02
+  vtl=0.0000000e+00 w0=0.0000000e+00 walpha0=-1.9557259e-13 wat=4.6564903e-01 wbeta0=5.3549638e-06
+  wint=2.1859000e-08 wk2=-9.2328587e-08 wketa=-9.0801561e-07 wkt1=-4.6564903e-07 wku0=0.0000000e+00
+  wkvth0=2.0000000e-07 wl=0.0000000e+00 wlc=0.0000000e+00 wln=1.0000000e+00 wlod=0.0000000e+00
+  wlodku0=1.0000000e+00 wlodvth=1.0000000e+00 wmax=1.2600000e-06 wmin=1.0000000e-06 wnfactor=-3.5019018e-05
+  wpclm=-5.0461019e-08 wr=1.0000000e+00 wu0=-2.5401808e-09 wua=2.5764227e-19 wub=1.1512823e-24
+  wuc=6.7910255e-16 wvsat=-4.6564499e-02 wvth0=5.3281370e-07 ww=0.0000000e+00 wwc=0.0000000e+00
+  wwl=0.0000000e+00 wwlc=0.0000000e+00 wwn=1.0000000e+00 xgl=0.0000000e+00 xgw=0.0000000e+00
+  xj=1.5000000e-07 xjbvs=1.0000000e+00 xl=0.0000000e+00 xn=3.0000000e+00 xpart=0.0000000e+00
+  xrcrg1=1.2000000e+01 xrcrg2=1.0000000e+00 xtis=2.0000000e+00 xw=0.0000000e+00

.model inverter:XM1:pfet_01v8:xsky130_fd_pr__pfet_01v8:sky130_fd_pr__pfet_01v8:msky130_fd_pr__pfet_01v8:sky130_fd_pr__pfet_01v8__model.62 pmos level=54 version=4.5 a0=-9.9544686e-01 a1=0.0000000e+00
+  a2=-3.9860003e+00 acde=8.0000000e-01 acnqsmod=0 af=1.0000000e+00 agidl=7.1279055e-09
+  ags=1.2500000e+00 aigbacc=4.3000000e-01 aigbinv=3.5000000e-01 aigc=4.3000000e-01 aigsd=4.3000000e-01
+  alpha0=1.0000000e-10 alpha1=1.0000000e-10 at=6.6598615e+05 b0=0.0000000e+00 b1=-4.6654513e-23
+  beta0=1.7668141e+01 bgidl=9.3461459e+08 bigbacc=5.4000000e-02 bigbinv=3.0000000e-02 bigc=5.4000000e-02
+  bigsd=5.4000000e-02 binunit=2 bvs=1.2690000e+01 capmod=2 cdsc=1.3000000e-04
+  cdscb=7.8000000e-04 cdscd=0.0000000e+00 cf=1.2000000e-11 cgbo=0.0000000e+00 cgdl=9.5482717e-12
+  cgdo=5.2489250e-11 cgidl=3.0000000e+02 cgsl=9.5482717e-12 cgso=5.2489250e-11 cigbacc=7.5000000e-02
+  cigbinv=6.0000000e-03 cigc=7.5000000e-02 cigsd=7.5000000e-02 cit=1.0000000e-05 cjs=7.3801945e-04
+  cjswgs=2.3915505e-10 cjsws=9.8888920e-11 ckappas=6.0000000e-01 clc=1.0000000e-07 cle=6.0000000e-01
+  delta=1.0000000e-02 diomod=1 dlc=-3.0000000e-09 dlcig=0.0000000e+00 dmcg=0.0000000e+00
+  dmcgt=0.0000000e+00 dmdg=0.0000000e+00 drout=1.0000000e+00 dsub=3.9026987e-01 dvt0=4.4955000e+00
+  dvt0w=-4.9772000e+00 dvt1=2.9400000e-01 dvt1w=1.1472000e+06 dvt2=1.5000000e-02 dvt2w=-8.9600000e-03
+  dvtp0=0.0000000e+00 dvtp1=0.0000000e+00 dwb=-1.7864000e-08 dwc=0.0000000e+00 dwg=-5.7220000e-09
+  ef=1.0000000e+00 egidl=1.0000000e-01 eigbinv=1.1000000e+00 em=4.1000000e+07 epsrox=3.9000000e+00
+  eta0=-2.8861269e+00 etab=-9.7918185e-01 eu=1.6700000e+00 fnoimod=1 fprout=0.0000000e+00
+  gbmin=1.0000000e-12 geomod=0 igbmod=0 igcmod=0 ijthsfwd=1.0000000e-01
+  ijthsrev=1.0000000e-01 jss=2.1483000e-05 jsws=8.0400000e-10 k1=-2.8786037e+00 k2=1.5858119e+00
+  k3=-1.5845000e+01 k3b=2.0000000e+00 keta=-9.8615600e-01 kf=0.0000000e+00 kt1=9.5239689e-01
+  kt1l=0.0000000e+00 kt2=-1.7698105e-01 ku0=4.5000000e-08 kvsat=5.0000000e-01 kvth0=3.2900000e-08
+  la0=2.6207616e-07 la2=9.5887991e-07 lagidl=-1.2859187e-15 lambda=0.0000000e+00 lat=-1.1821557e-01
+  lb1=8.3039435e-30 lbeta0=-2.0307064e-06 lbgidl=1.1637818e+01 lc=5.0000000e-09 ldsub=-2.3186474e-08
+  leta0=6.1863802e-07 letab=1.5627874e-07 lint=-1.3994000e-08 lintnoi=-2.0000000e-07 lk1=7.5411139e-07
+  lk2=-3.4521058e-07 lketa=2.0793478e-07 lkt1=-2.9584398e-07 lkt2=1.0141942e-08 lku0=0.0000000e+00
+  lkvth0=0.0000000e+00 ll=0.0000000e+00 llc=0.0000000e+00 lln=1.0000000e+00 llodku0=0.0000000e+00
+  llodvth=0.0000000e+00 lmax=1.8000000e-07 lmin=1.5000000e-07 lnfactor=8.0282415e-07 lodeta0=1.0000000e+00
+  lodk2=1.0000000e+00 lp=1.0000000e+00 lpclm=-7.5813905e-07 lpdiblc1=-7.9488155e-07 lpdiblc2=-1.9935289e-08
+  lpdiblcb=3.0385009e-07 lpe0=0.0000000e+00 lpeb=0.0000000e+00 lpscbe2=2.7340905e-17 lu0=-2.6081666e-09
+  lua=-9.8182197e-16 lua1=2.7619141e-17 lub=9.9860379e-25 lub1=1.5308793e-25 luc=-5.6460284e-19
+  luc1=8.5595572e-18 lute=4.3842950e-07 lvoff=-3.7058686e-08 lvsat=-1.1496936e-01 lvth0=9.2039115e-08
+  lw=0.0000000e+00 lwc=0.0000000e+00 lwl=0.0000000e+00 lwlc=0.0000000e+00 lwn=1.0000000e+00
+  minv=0.0000000e+00 mjs=3.4629000e-01 mjswgs=9.2740000e-01 mjsws=2.9781000e-01 mobmod=0
+  moin=1.8130000e+01 ndep=1.7000000e+17 nfactor=-2.5202305e+00 ngate=1.0000000e+23 ngcon=1.0000000e+00
+  nigbacc=1.0000000e+00 nigbinv=3.0000000e+00 nigc=1.0000000e+00 njs=1.3632000e+00 noff=3.9000000e+00
+  noia=1.5000000e+42 noib=0.0000000e+00 noic=0.0000000e+00 nsd=1.0000000e+20 ntnoi=1.0000000e+00
+  ntox=1.0000000e+00 pa0=-5.9401795e-13 pa2=-9.0698822e-13 pagidl=2.0637229e-21 pat=1.3462002e-07
+  pb1=-1.3580204e-35 pbeta0=1.2162406e-12 pbgidl=-1.9032396e-05 pbs=6.5870000e-01 pbswgs=1.4338000e+00
+  pbsws=7.4180000e-01 pclm=4.3041982e+00 pdiblc1=4.0937644e+00 pdiblc2=1.0534151e-01 pdiblcb=-1.2222147e+00
+  pdits=0.0000000e+00 pditsd=0.0000000e+00 pditsl=0.0000000e+00 pdsub=1.4296272e-14 permod=1
+  peta0=-7.7155733e-13 petab=-1.6877001e-13 phin=0.0000000e+00 pigcd=1.0000000e+00 pk1=-6.5240830e-13
+  pk2=3.1846147e-13 pketa=-3.3209256e-13 pkt1=2.5828484e-13 pkt2=-1.2630696e-14 pku0=0.0000000e+00
+  pkvth0=0.0000000e+00 pnfactor=-6.2606879e-13 poxedge=1.0000000e+00 ppclm=9.3533260e-13 ppdiblc1=9.7443098e-13
+  ppdiblc2=2.5343649e-14 ppdiblcb=-4.9657258e-13 ppscbe2=-3.5606189e-22 prt=0.0000000e+00 prwb=-3.2348000e-01
+  prwg=1.3760000e-01 pscbe1=8.0000000e+08 pscbe2=9.6284831e-09 pu0=3.1656648e-15 pua=1.1048237e-21
+  pua1=1.5595043e-23 pub=-1.0498151e-30 pub1=-2.9836797e-31 puc=5.9895453e-25 puc1=-2.1968389e-24
+  pute=-5.4028446e-13 pvag=0.0000000e+00 pvoff=4.5217955e-14 pvsat=1.1716259e-07 pvth0=-1.6870743e-13
+  rbdb=5.0000000e+01 rbodymod=1 rbpb=5.0000000e+01 rbpd=5.0000000e+01 rbps=5.0000000e+01
+  rbsb=5.0000000e+01 rdsmod=0 rdsw=5.4788000e+02 rdswmin=0.0000000e+00 rdw=0.0000000e+00
+  rdwmin=0.0000000e+00 rgatemod=0 rnoia=6.9000000e-01 rnoib=3.4000000e-01 rsh=1.0000000e+00
+  rshg=1.0000000e-01 rsw=0.0000000e+00 rswmin=0.0000000e+00 saref=1.0400000e-06 sbref=1.0400000e-06
+  steta0=0.0000000e+00 stk2=0.0000000e+00 tcj=1.2407000e-03 tcjsw=3.7357000e-04 tcjswg=2.0000000e-12
+  tempmod=0 tku0=0.0000000e+00 tnoia=2.5000000e+07 tnoib=0.0000000e+00 tnoimod=1
+  tnom=3.0000000e+01 toxe=4.2300000e-09 toxm=4.2300000e-09 toxref=4.2300000e-09 tpb=2.0386000e-03
+  tpbsw=1.2460000e-03 tpbswg=0.0000000e+00 trnqsmod=0 tvfbsdoff=0.0000000e+00 tvoff=0.0000000e+00
+  u0=1.7981468e-02 ua=2.9137552e-09 ua1=-4.8881808e-11 ub=-3.1786562e-18 ub1=-4.9119253e-19
+  uc=3.0410342e-12 uc1=-4.1642242e-11 ud=0.0000000e+00 up=0.0000000e+00 ute=-2.6756831e+00
+  vbm=-3.0000000e+00 vfbcv=-1.4469000e-01 vfbsdoff=0.0000000e+00 voff=-1.0975886e-01 voffcv=-1.0701000e-01
+  voffl=0.0000000e+00 vsat=6.3398740e+05 vth0=-1.5022826e+00 vtl=0.0000000e+00 w0=0.0000000e+00
+  wa0=3.8802216e-06 wa2=4.4386354e-06 wagidl=-1.0974982e-14 wat=-6.9515330e-01 wb1=7.6298427e-29
+  wbeta0=-4.7419822e-06 wbgidl=1.0693078e+02 wdsub=-8.0321550e-08 weta0=3.8629364e-06 wetab=1.0558414e-06
+  wint=7.3039000e-09 wk1=3.6118907e-06 wk2=-1.7191698e-06 wketa=1.6135470e-06 wkt1=-1.4511363e-06
+  wkt2=7.0963749e-08 wku0=2.5000000e-07 wkvth0=2.0000000e-07 wl=0.0000000e+00 wlc=0.0000000e+00
+  wln=1.0000000e+00 wlod=0.0000000e+00 wlodku0=1.0000000e+00 wlodvth=1.0000000e+00 wmax=1.6500000e-06
+  wmin=1.2600000e-06 wnfactor=4.2279219e-06 wpclm=-4.5431672e-06 wpdiblc1=-4.8341773e-06 wpdiblc2=-1.3079138e-07
+  wpdiblcb=1.9968422e-06 wpscbe2=1.2491480e-15 wr=1.0000000e+00 wu0=-1.8314488e-08 wua=-6.0206570e-15
+  wua1=7.9499443e-18 wub=5.7434823e-24 wub1=1.6763375e-24 wuc=-3.0009336e-18 wuc1=1.2342624e-17
+  wute=3.0355106e-06 wvoff=-3.1479708e-07 wvsat=-5.3746632e-01 wvth0=8.9297031e-07 ww=0.0000000e+00
+  wwc=0.0000000e+00 wwl=0.0000000e+00 wwlc=0.0000000e+00 wwn=1.0000000e+00 xgl=0.0000000e+00
+  xgw=0.0000000e+00 xj=1.5000000e-07 xjbvs=1.0000000e+00 xl=0.0000000e+00 xn=3.0000000e+00
+  xpart=0.0000000e+00 xrcrg1=1.2000000e+01 xrcrg2=1.0000000e+00 xtis=5.2000000e+00 xw=0.0000000e+00

* end of model section

.option autostop numdgt=6 measdgt=6 ingold=2 save=nooutput
.tran 1.00e-12 1.0000000e-10 

.end

* end of sim.sp
